module test(





);
endmodule